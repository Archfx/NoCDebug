// megafunction wizard: %Virtual JTAG%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: sld_virtual_jtag 

// ============================================================
// File Name: vjtag.v
// Megafunction Name(s):
// 			sld_virtual_jtag
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 13.0.0 Build 156 04/24/2013 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2013 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.





module vjtag #(
	parameter  VJTAG_INDEX=126

)(
	ir_out,
	tdo,
	ir_in,
	tck,
	tdi,
	virtual_state_cdr,
	virtual_state_cir,
	virtual_state_e1dr,
	virtual_state_e2dr,
	virtual_state_pdr,
	virtual_state_sdr,
	virtual_state_udr,
	virtual_state_uir);

	input	[2:0]  ir_out;
	input	  tdo;
	output	[2:0]  ir_in;
	output	  tck;
	output	  tdi;
	output	  virtual_state_cdr;
	output	  virtual_state_cir;
	output	  virtual_state_e1dr;
	output	  virtual_state_e2dr;
	output	  virtual_state_pdr;
	output	  virtual_state_sdr;
	output	  virtual_state_udr;
	output	  virtual_state_uir;

	wire  sub_wire0;
	wire  sub_wire1;
	wire [2:0] sub_wire2;
	wire  sub_wire3;
	wire  sub_wire4;
	wire  sub_wire5;
	wire  sub_wire6;
	wire  sub_wire7;
	wire  sub_wire8;
	wire  sub_wire9;
	wire  sub_wire10;
	wire  virtual_state_cir = sub_wire0;
	wire  virtual_state_pdr = sub_wire1;
	wire [2:0] ir_in = sub_wire2[2:0];
	wire  tdi = sub_wire3;
	wire  virtual_state_udr = sub_wire4;
	wire  tck = sub_wire5;
	wire  virtual_state_e1dr = sub_wire6;
	wire  virtual_state_uir = sub_wire7;
	wire  virtual_state_cdr = sub_wire8;
	wire  virtual_state_e2dr = sub_wire9;
	wire  virtual_state_sdr = sub_wire10;

// `ifndef VERILATOR
// `ifndef MODEL_TECH
// 	// sld_virtual_jtag	sld_virtual_jtag_component (
// 	// 			.ir_out (ir_out),
// 	// 			.tdo (tdo),
// 	// 			.virtual_state_cir (sub_wire0),
// 	// 			.virtual_state_pdr (sub_wire1),
// 	// 			.ir_in (sub_wire2),
// 	// 			.tdi (sub_wire3),
// 	// 			.virtual_state_udr (sub_wire4),
// 	// 			.tck (sub_wire5),
// 	// 			.virtual_state_e1dr (sub_wire6),
// 	// 			.virtual_state_uir (sub_wire7),
// 	// 			.virtual_state_cdr (sub_wire8),
// 	// 			.virtual_state_e2dr (sub_wire9),
// 	// 			.virtual_state_sdr (sub_wire10)
// 	// 			);


// 	defparam
// 		sld_virtual_jtag_component.sld_auto_instance_index = "NO",
// 		sld_virtual_jtag_component.sld_instance_index = VJTAG_INDEX,
// 		sld_virtual_jtag_component.sld_ir_width = 3,
// 		sld_virtual_jtag_component.sld_sim_action = "((0,1,7,3),(0,2,ff,20),(0,1,6,3),(0,2,ffffffff,20),(0,2,1,20),(0,2,2,20),(0,2,3,20),(0,2,4,20))",
// 		sld_virtual_jtag_component.sld_sim_n_scan = 8,
// 		sld_virtual_jtag_component.sld_sim_total_length = 198;
// `endif //MODEL_TECH
// `endif //VERILATOR

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
// Retrieval info: PRIVATE: show_jtag_state STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: SLD_AUTO_INSTANCE_INDEX STRING "NO"
// Retrieval info: CONSTANT: SLD_INSTANCE_INDEX NUMERIC "126"
// Retrieval info: CONSTANT: SLD_IR_WIDTH NUMERIC "3"
// Retrieval info: CONSTANT: SLD_SIM_ACTION STRING "((0,1,7,3),(0,2,ff,20),(0,1,6,3),(0,2,ffffffff,20),(0,2,1,20),(0,2,2,20),(0,2,3,20),(0,2,4,20))"
// Retrieval info: CONSTANT: SLD_SIM_N_SCAN NUMERIC "8"
// Retrieval info: CONSTANT: SLD_SIM_TOTAL_LENGTH NUMERIC "198"
// Retrieval info: USED_PORT: ir_in 0 0 3 0 OUTPUT NODEFVAL "ir_in[2..0]"
// Retrieval info: USED_PORT: ir_out 0 0 3 0 INPUT NODEFVAL "ir_out[2..0]"
// Retrieval info: USED_PORT: tck 0 0 0 0 OUTPUT NODEFVAL "tck"
// Retrieval info: USED_PORT: tdi 0 0 0 0 OUTPUT NODEFVAL "tdi"
// Retrieval info: USED_PORT: tdo 0 0 0 0 INPUT NODEFVAL "tdo"
// Retrieval info: USED_PORT: virtual_state_cdr 0 0 0 0 OUTPUT NODEFVAL "virtual_state_cdr"
// Retrieval info: USED_PORT: virtual_state_cir 0 0 0 0 OUTPUT NODEFVAL "virtual_state_cir"
// Retrieval info: USED_PORT: virtual_state_e1dr 0 0 0 0 OUTPUT NODEFVAL "virtual_state_e1dr"
// Retrieval info: USED_PORT: virtual_state_e2dr 0 0 0 0 OUTPUT NODEFVAL "virtual_state_e2dr"
// Retrieval info: USED_PORT: virtual_state_pdr 0 0 0 0 OUTPUT NODEFVAL "virtual_state_pdr"
// Retrieval info: USED_PORT: virtual_state_sdr 0 0 0 0 OUTPUT NODEFVAL "virtual_state_sdr"
// Retrieval info: USED_PORT: virtual_state_udr 0 0 0 0 OUTPUT NODEFVAL "virtual_state_udr"
// Retrieval info: USED_PORT: virtual_state_uir 0 0 0 0 OUTPUT NODEFVAL "virtual_state_uir"
// Retrieval info: CONNECT: @ir_out 0 0 3 0 ir_out 0 0 3 0
// Retrieval info: CONNECT: @tdo 0 0 0 0 tdo 0 0 0 0
// Retrieval info: CONNECT: ir_in 0 0 3 0 @ir_in 0 0 3 0
// Retrieval info: CONNECT: tck 0 0 0 0 @tck 0 0 0 0
// Retrieval info: CONNECT: tdi 0 0 0 0 @tdi 0 0 0 0
// Retrieval info: CONNECT: virtual_state_cdr 0 0 0 0 @virtual_state_cdr 0 0 0 0
// Retrieval info: CONNECT: virtual_state_cir 0 0 0 0 @virtual_state_cir 0 0 0 0
// Retrieval info: CONNECT: virtual_state_e1dr 0 0 0 0 @virtual_state_e1dr 0 0 0 0
// Retrieval info: CONNECT: virtual_state_e2dr 0 0 0 0 @virtual_state_e2dr 0 0 0 0
// Retrieval info: CONNECT: virtual_state_pdr 0 0 0 0 @virtual_state_pdr 0 0 0 0
// Retrieval info: CONNECT: virtual_state_sdr 0 0 0 0 @virtual_state_sdr 0 0 0 0
// Retrieval info: CONNECT: virtual_state_udr 0 0 0 0 @virtual_state_udr 0 0 0 0
// Retrieval info: CONNECT: virtual_state_uir 0 0 0 0 @virtual_state_uir 0 0 0 0
// Retrieval info: GEN_FILE: TYPE_NORMAL vjtag.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL vjtag.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL vjtag.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL vjtag.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL vjtag_inst.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL vjtag_bb.v TRUE
// Retrieval info: LIB_FILE: altera_mf
